netcdf sofa {
		// This is a SOFA file
:Conventions="SOFA";

		// global attributes
:SOFAConvention="SimpleFreeFieldHRTF";
:SOFAConventionVersion="0.0.1";
:ApplicationName="ncgen";
:ApplicationVersion="0.0.0";
:AuthorContact="piotr@majdak.com";
:Licence="CC BY-SA 3.0";
:Organization="ARI, OeAW";
:DatabaseName="ARI";
:SubjectID="template";

dimensions: 
N = unlimited, M=unlimited; C=3;	// SOFA defined
R=2, E=1; // Measurement specific

variables:
		// general dimensions
int		R(R),E(E),M(M),C(C),N(N);
R:LongName="number of receivers";
E:LongName="number of emitters";
M:LongName="number of measurements";
C:LongName="coordinate triplet";

		// Data-type
:DataType="FIR";
float	Data.IR(M,R,N);
float	Data.SamplingRate;
N:LongName="time";
N:Units="samples";
Data.SamplingRate:Units="hertz";

		// Listener
float	ListenerPosition(M,C);
ListenerPosition:Type="cartesian";
ListenerPosition:Units="meter";
float	ListenerUp(M,C);
ListenerUp:Type="cartesian";
ListenerUp:Units="meter";
float	ListenerView(M,C);
ListenerView:Type="cartesian";
ListenerView:Units="meter";
float	ListenerRotation(M,C);
ListenerRotation:Type="din9300";
ListenerPosition:Type="degrees";

		// Receivers
float	ReceiverPosition(R,C);
ReceiverPosition:Type="cartesian";
ReceiverPosition:Units="meter";

		// Source
float	SourcePosition(C);
SourcePosition:Type="cartesian";
SourcePosition:Units="meter";
float	SourceUp(C);
SourceUp:Type="cartesian";
SourceUp:Units="meter";
float	SourceView(C);
SourceView:Type="cartesian";
SourceView:Units="meter";

		// Emitters
float 	EmitterPosition(C);
EmitterPosition:Type="cartesian";
EmitterPosition:Units="meter";

		// Room
:RoomType="free field";
		
data:
	SourcePosition=0,0,0;
	SourceUp=0,0,1;
	SourceView=1,0,0;
	EmitterPosition=0,0,0;
	ListenerPosition=1.2,0,0;
	ListenerView=0,0,0;
	ListenerUp=1.2,0,0;
	ReceiverPosition=0,-0.09,0 ,0,0.09,0;
}
